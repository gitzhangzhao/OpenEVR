--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:    09:11:20 10/18/05
-- Design Name:    
-- Module Name:    gtl_all - Behavioral
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity vmesimple is
port
(
    -- System clock input : 50MHz clock used
   clk_i                         :  in    std_logic;
    -- VME signals
	DATA									:	inout		std_logic_vector(31 downto 0);
	BERR									:	out		std_logic;
	DTACK									:	out		std_logic;
	ADDR									:	in			std_logic_vector(23 downto 1);
	WRITE2_BAR							:	in			std_logic;
	AM_LV									:	in			std_logic_vector(5 downto 0);
	IACKIN_BAR							:	in			std_logic;
	IACK_BAR								:	in			std_logic;
	GA_LV									:	in			std_logic_vector(4 downto 0);
	DS0_BAR								:	in			std_logic;
	DS1_BAR								:	in			std_logic;
	LWORD_BAR							:	in			std_logic;
	SYSRESET_BAR						:	in			std_logic;
	AS_BAR								:	in			std_logic;
	IACKOUT_BAR							:	out		std_logic;
    -- VME signals end here

    -- VME buffers
   VME_DTACK_OE_o  : out std_logic;
   VME_DATA_DIR_o  : out std_logic;
   VME_DATA_OE_N_o : out std_logic;
   VME_ADDR_DIR_o  : out std_logic;
   VME_ADDR_OE_N_o : out std_logic;
	
	--VME module output signals of register set
	addr_dma1_o		 : out std_logic_vector(18 downto 2);
	--register02_addr : out std_logic_vector(18 downto 2);
	data_wr_o       : out std_logic_vector(31 downto 0);
	data_rd_i		 : in  std_logic_vector(31 downto 0);
	--write_int_o		: out std_logic;
	ds_dly_clk_o    : out std_logic;
	board_sel_o		 : out std_logic
	
	--VME module output signals of mappingRAM
	--mappingRAM_board_sel		:   out std_logic
	 
	);	
end vmesimple;

architecture Behavioral of vmesimple is

	attribute BOX_TYPE   : STRING ;
   component BUFG
      port ( I : in    std_logic; 
             O : out   std_logic);
   end component;
   attribute BOX_TYPE of BUFG : COMPONENT is "BLACK_BOX";
   
   
   component IO32_PORTS
   port(I   : in    std_logic_vector(31 downto 0);
	     O   : out   std_logic_vector(31 downto 0);
		  T   : in    std_logic;
		  IO  : inout std_logic_vector(31 downto 0)
		  );
  end component;
	
	
	
-- Global clock buffered by bufg
	signal	CLK_Global						:	std_logic;
	
	-- VME related signals
	--signal data_wr, data_rd					:			std_logic_vector(15 downto 0);
	signal data_bus_read_ena_bar			:			std_logic;
	signal addr_reg							:			std_logic_vector(23 downto 0);
	signal addr_dma1							:			std_logic_vector(18 downto 2);
	signal cnt_addr_dma						:			std_logic_vector(16 downto 0);
	signal as_int								:			std_logic;
	signal AM_LV_reg							:			std_logic_vector(5 downto 0);
	signal GA_LV_int							:			std_logic_vector(4 downto 0);
	signal write_int							:			std_logic;
	signal ds0_int								:			std_logic;
	signal ds1_int								:			std_logic;
	signal ds_int								:			std_logic;
	signal ds_dly1								:			std_logic;
	signal ds_dly2								:			std_logic;
	signal ds_dly3								:			std_logic;
	signal ds_dly4								:			std_logic;
	signal ds_dly5								:			std_logic;
	signal ds_dly6								:			std_logic;
	signal ds_dly7								:			std_logic;
	signal ds_dly8								:			std_logic;
	signal ds_dly9								:			std_logic;
	signal ds_dly10							:			std_logic;
	signal ds_dly_clk							:			std_logic;
	signal board_sel							:			std_logic;
	signal dtack_int							:			std_logic;
	-- reset signal generated by VME operation	
	signal reset_vme							:			std_logic;
	-- VME related signals end here


begin
    
    VME_ADDR_DIR_o  <= '0';
    VME_ADDR_OE_N_o <= '0';
	 
	 addr_dma1_o     <= addr_dma1;
	 --data_wr_o       <= data_wr;
	 --data_rd         <= data_rd_i;
	 --write_int_o     <= write_int;
	 ds_dly_clk_o    <= ds_dly_clk;
	 board_sel_o     <= board_sel;


-- clock fanout
	clock_buffer : bufg
   port map(i  => clk_i
	        ,o  => CLK_Global
			  );
	
-- VME operations
	-- data ports mapping
	data_bus_read_ena_bar <= not (board_sel and (not write_int));

	DATA_BUS32_IOs : IO32_PORTS
   port map(I  => data_rd_i
	        ,O  => data_wr_o
			  ,IO => data
			  ,T  => data_bus_read_ena_bar
			  );
	-- data ports mapping end here

	-- AS registered by internal clock
	AS_register_generation : process(AS_BAR, CLK_Global)
	begin
		if(CLK_Global'event and CLK_Global = '1') then
			as_int	<= not AS_BAR;
		end if;
	end process;	
	-- -- --

	-- write signal 
	write_int <= not WRITE2_BAR;
	-- write signal end here
	
	-- DS registered by internal clock
	DS_register_generation : process(DS0_BAR, DS1_BAR, CLK_Global)
	begin
		if(CLK_Global'event and CLK_Global = '1') then
			ds0_int	<= not DS0_BAR;
			ds1_int	<= not DS1_BAR;
		end if;
	end process;	

	ds_int	<= ds0_int and ds1_int;

	ds_internal_delay : process(CLK_Global)
	begin
		if(CLK_Global'event and CLK_Global = '1') then
			ds_dly1		<= ds_int;
			ds_dly2		<= ds_dly1;
			ds_dly3		<= ds_dly2;
			ds_dly4		<= ds_dly3;
			ds_dly5		<= ds_dly4;
			ds_dly6		<= ds_dly5;
			ds_dly7		<= ds_dly6;
			ds_dly8		<= ds_dly7;
			ds_dly9		<= ds_dly8;
			ds_dly10		<= ds_dly9;
		end if;
	end process;
	
	ds_dly_clk	<= ds_dly3;
	
	-- -- --
	
	-- dtack generation from here
	dtack <= not dtack_int;
	VME_DTACK_OE_o <= not board_sel;

	dtack_internal_generation : process(ds_dly6, board_sel, ds_int) 
	begin
		if(ds_int = '0') then
			dtack_int <= '0';
		else
			if(board_sel = '1') then
				if(ds_dly6'event and ds_dly6 = '1') then
					dtack_int <= '1';
				end if;
			end if;
		end if;
	end process;
	-- dtack generation end here
	
	-- ADDR registered by as_int
	addr_register_generation : process(as_int, ADDR, LWORD_BAR, AM_LV)
	begin
		if(as_int'event and as_int = '1') then
			addr_reg(23 downto 1)	<= addr;
			addr_reg(0)					<= LWORD_BAR;
			AM_LV_reg					<= AM_LV;
		end if;
	end process;	
	-- -- --

	-- Board Gates -- [4 : 0] corresponding to Addr [23 : 19]
	GA_LV_int(0)	<= not GA_LV(0);
	GA_LV_int(1)	<= not GA_LV(1);
	GA_LV_int(2)	<= not GA_LV(2);
	GA_LV_int(3)	<= not GA_LV(3);
	--GA_LV_int(4)	<= not GA_LV(4);
	--GA_LV_int(0)	<= '1';
	--GA_LV_int(1)	<= '1';
	--GA_LV_int(2)	<= '0';
	--GA_LV_int(3)	<= '0';
	GA_LV_int(4)	<= '0';
--	-- -- --

	-- Board selection determination
	board_selection_judge : process(addr_reg, GA_LV_int, AM_LV_reg)
	begin
		if((addr_reg(23 downto 19) = GA_LV_int) and (addr_reg(1 downto 0) = "00") and
												(AM_LV_reg >= "111000" and AM_LV_reg <= "111111")) then
			board_sel	<= '1';
		else
			board_sel	<= '0';
		end if;
	end process;
	
	
	--BS_BAR	<= not board_sel;
	VME_DATA_OE_N_o <= not board_sel;
	VME_DATA_DIR_o  <= WRITE2_BAR;
	-- -- --

	-- DMA address generation
	addr_dma1	     <=	addr_reg(18 downto 2) + cnt_addr_dma;
	--register02_addr  <=	addr_reg(18 downto 2);

	DMA_address_generation_add : process(as_int, dtack_int)
	begin
		if(as_int = '0') then
			cnt_addr_dma <= (others => '0');
		else
			if(dtack_int'event and dtack_int = '0') then
				cnt_addr_dma	<= cnt_addr_dma + 1;
			end if;
		end if;
	end process;
	-- -- --

	VME_reset_generation : process(CLK_Global, board_sel, write_int, ds_dly_clk, addr_dma1)
	begin
		if(CLK_Global'event and CLK_Global = '1') then
			if(addr_dma1 = '1' & X"ffff") then
				reset_vme <= board_sel and write_int and ds_dly_clk;
			else
				reset_vme <= '0';
			end if;
		end if;
	end process;
	

--mappingRAM selection judge
--   mappingRAM_board_selection_judge : process(addr_dma1, board_sel)
--	begin
--      if (addr_dma1 > '0' & X"000f" and addr_dma1 < '0'& X"010f" and board_sel = '1') then
--          mappingRAM_board_sel <= '1';
--		else
--		    mappingRAM_board_sel <= '0';
--		end if;
--	end process;
	
	
	-- bus interrupt related from here
	IACKOUT_BAR <= IACKIN_BAR;
	--IRQ_Board	<= '0';
	BERR			<= '1';
	-- bus interrupt related end here

-- VME operations end here



end Behavioral;

